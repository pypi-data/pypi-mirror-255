netcdf base {

dimensions:
	time = UNLIMITED ; # Main dimension

variables:

	string station_name;
	    station_name:standard_name = "platform_name" ;
		station_name:long_name = "station_name" ;
		station_name:cf_role = "timeseries_id" ;

    float latitude ;
		latitude:long_name = "station latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:_CoordinateAxisType = "Lat" ;
		latitude:axis = "Y" ;

	float longitude ;
		longitude:long_name = "station longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:_CoordinateAxisType = "Lon" ;
		longitude:axis = "X" ;

	float elevation;
		elevation:long_name = "Elevation above mean seal level" ;
		elevation:standard_name = "height_above_mean_sea_level" ;
		elevation:units = "m" ;
		elevation:axis = "Z" ;

	double crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = "0.0" ;
		crs:semi_major_axis = "6378137.0" ;
		crs:inverse_flattening = "298.257223563" ;
		crs:epsg_code = "EPSG:4326";

	uint Time(time) ;
		Time:long_name = "Time of measurement" ;
		Time:standard_name = "time" ;
		Time:units = "seconds since 1970-01-01 00:00:00";
		Time:time_origin = "1970-01-01 00:00:00" ;
		Time:time_zone= "UTC"
		Time:abbreviation = "Date/Time" ;
		Time:axis = "T" ;
		Time:calendar = "gregorian" ;

    float GHI(time) ;
		GHI:long_name = "Global Horizontal Irradiance" ;
		GHI:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		GHI:abbreviation = "SWD" ;
		GHI:units = "W m-2" ;
		GHI:_valid_min=0.0 ;
		GHI:_valid_max=3000 ;
		GHI:grid_mapping = "crs" ;
		GHI:least_significant_digit=1;

	float DIF(time) ;
		DIF:long_name = "Diffuse horizontal radiation" ;
		DIF:standard_name = "surface_diffuse_downwelling_shortwave_flux_in_air" ;
		DIF:abbreviation = "DHI" ;
		DIF:units = "W m-2" ;
		DIF:_valid_min=0.0 ;
		DIF:_valid_max=3000 ;
		DIF:grid_mapping = "crs" ;
		DIF:least_significant_digit=1;

	float DNI(time) ;
		DNI:long_name = "Beam (or direct) normal radiation" ;
		DNI:standard_name = "direct_downwelling_shortwave_flux_in_air" ;
		DNI:abbreviation = "BNI" ;
		DNI:units = "W m-2" ;
		DNI:_valid_min=0.0 ;
		DNI:_valid_max=3000 ;
		DNI:grid_mapping = "crs" ;
		DNI:least_significant_digit=1;

	float GHIcalc(time) ;
		GHIcalc:parameter = "Short-wave downward (GLOBAL) radiation" ;
		GHIcalc:long_name = "Global Horizontal Irradiance calculated with the diffuse and direct components" ;
		GHIcalc:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		GHIcalc:abbreviation = "SWD" ;
		GHIcalc:units = "W m-2" ;
		GHIcalc:_valid_min = -10. ;
		GHIcalc:_valid_max = 3000 ;
		GHIcalc:least_significant_digit = 1 ;

    float Elev(time) ;
		Elev:parameter = "Solar elevation angle" ;
		Elev:long_name = "Solar elevation angle" ;
		Elev:abbreviation = "Elev" ;
		Elev:units = "degree" ;
		Elev:_valid_min = -1 ;
		Elev:_valid_max = 95 ;
		Elev:least_significant_digit = 3 ;

	float Azim(time) ;
		Azim:parameter = "Solar azimuth angle" ;
		Azim:long_name = "Solar azimuth angle" ;
		Azim:abbreviation = "Azim" ;
		Azim:units = "degree" ;
		Azim:_valid_min = -362 ;
		Azim:_valid_max = 362 ;
		Azim:least_significant_digit = 3 ;

	float Kc(time) ;
		Kc:parameter = "Clear sky index" ;
		Kc:long_name = "Clear sky index" ;
		Kc:abbreviation = "Kc" ;
		Kc:comment = "Kc is the clearsky index calculated with CAMS mcclear with GHIcalc/GHI McClear" ;
		Kc:_valid_min = -0.1 ;
		Kc:_valid_max = 2 ;
		Kc:least_significant_digit = 3 ;
		
	int flagPPLDIF(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;
		
	int flagERLDIF(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagPPLDNI(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagERLDNI(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagPPLGHI(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagERLGHI(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flag3highSZA(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flag3lowSZA(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKt(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKKt(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKn(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKnKt(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKhighSZA(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagKlowSZA(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagTracker(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;

	int flagManual(time) ;
		*:_valid_min =  0;
		*:_valid_max =  1;
		*:_FillValue = -999;
		*:missing_value = -999;



# Global attributes

    # Main info
    :id = "{Network_ID}-{Station_ID}";
    :title = "Timeseries of {Network_LongName} ({Network_ID}). Station : {Station_Name}" ;
    :description = "Reference data used for the validation work in the IEA PVPS task 16" ;
    :featureType = "timeSeries" ;
    :cdm_data_type = "timeSeries";

    # Conventions
    :Conventions = "CF-1.9,ACDD-1.3";

    # Publisher [ACDD1.3]
    :publisher_name = "Lionel MENARD, Raphael JOLIVET, Yves-Marie SAINT-DRENAN, Philippe BLANC";
    :publisher_email = "lionel.menard@mines-paristech.fr, raphael.jolivet@mines-paristech.fr, saint-drenan@mines-paristech.fr, philippe.blanc@mines-paristech.fr";
    :publisher_url = "https://www.oie.minesparis.psl.eu/" ;
    :publisher_institution = "Mines Paristech - PSL"

    # Creator info [ACDD1.3]
    :creator_name =  "{Station_ContactName}" ;
    :institution =  "{Station_Institute}" ;
    :metadata_link =  "{Station_Url}";
    :creator_url = "{Network_DescriptionURL}" ;
    :creator_email = "{Network_ContactPersonMail}";
    :references = "{Network_References}" ;
    :license = "{Network_LicenseInfoURL}" ;

    :comment = "{Station_Comment}" ;

    # Station info & coordinates [ACDD1.3]
    :project = "IEA PVPS task 16"; # Network long name
    :platform = "{Station_Name}" ; # Should be a long / full name
    :geospatial_lat_min = {Station_Latitude} ;
    :geospatial_lon_min = {Station_Longitude} ;
    :geospatial_lat_max = {Station_Latitude} ;
    :geospatial_lon_max = {Station_Longitude} ;
    :geospatial_vertical_min = {Station_Elevation};
    :geospatial_vertical_max = {Station_Elevation};
    :geospatial_bounds = "POINT({Station_Latitude} {Station_Longitude})";
    :geospatial_bounds_crs = "EPSG:4326";

    # Time information
    :time_coverage_start = "{Station_StartDate}T00:00:00" ;  # First data [Dataset Discovery v1.0]
    :time_coverage_end = "{Station_EndDate}T00:00:00";  # Last data [Dataset Discovery v1.0]
    :time_coverage_resolution = "P{Station_TimeResolution}"; # Resolution in  ISO 8601:2004 duration format [Dataset Discovery v1.0]
    :local_time_zone = "{Station_Timezone}" ;
    :date_created = "{CreationTime}";
    :date_modified = "{UpdateTime}";

    #
    # -- Additional metadata (custom to insitu)
    #

    # IDs
    :network_id = "{Network_ID}"; # Short ID
    :station_id = "{Station_ID}"; # Short ID
    :station_uid = "{Station_UID}" ; # Numeric ID, if any
    :station_wmo_id =  "{Station_WMOID}"; # WMO ID, if any

    # Surface
    :surface_type = "{Station_SurfaceType}" ; # rock, gress, concrete, cultivated, ...
    :topography_type = "{Station_TopographyType}" ; # flat, hilly, moutain valley, mountain top, ...
    :rural_urban = "{Station_RuralUrban}" ; # "rural" or "urban"

    # Location of station
    :network_region = "{Network_Region}";
    :station_address =  "{Station_Address}" ;
    :station_city =  "{Station_City}" ;
    :station_country =  "{Station_Country}" ;

    # Commission / decommission dates
    :station_commision_date  =  "{Station_CommissionDate}";
    :station_decommision_date =  "{Station_DecommissionDate}";

    # Misc
    :climate = "{Station_Climate}" ; # KoeppenGeiger climate at location of the station
    :operation_status =  "{Station_OperationStatus}";



}
